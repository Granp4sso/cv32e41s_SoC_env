// Copyright 2023 University of Naples, Federico II
// Date: 09 October 2023

////////////////////////////////////////////////////////////////////////////////
//                                                                            //
// Engineer:       Stefano Mercogliano - stefano.mercogliano@unina.it         //
//                                                                            //
//                                                                            //
// Description:    SPI Slave Interface                                        //        
//                                                                            //
////////////////////////////////////////////////////////////////////////////////